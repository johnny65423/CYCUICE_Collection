
module And(a, b, out);

    input a, b;
    output out;

    and(out,a,b);

endmodule

