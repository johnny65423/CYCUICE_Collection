
module Or(a, b, out);

    input a, b;
    output out;
   
    or(out,a,b);

endmodule
